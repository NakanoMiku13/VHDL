library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity ROM is
	Port(
		direction : in std_logic_vector(4 downto 0);
		memoryValue : out std_logic_vector(28 downto 0)
	);
end ROM;
architecture ArchROM of ROM is
	type Rom_instrucciones is array(0 to 31) of std_logic_vector(28 downto 0);
	constant TR : Rom_instrucciones := (
	--Instrucciones tipo R
		0  => "00000000000000000000000000000",
		1  => "00000101000100010000000000000",
		2  => "00001010001000100000000000000",
		3  => "00001111001100110000000000000",
		4  => "00010000010001000000000000000",
		5  => "00010100100101010000000000000",
		6  => "00011000111001100000000000000",
		7  => "00011111111101110000000000000",
		8  => "00100011100010000000000000000",
		9  => "00100111010110010000000000000",
		--Instruccines tipo I
		10 => "00101001010110000000000000000",
		11 => "00101110100111000000000000000",
		12 => "00110011111000000000000000000",
		--Instruccines tipo J
		13 => "00110100010000000000000000000",
		14 => "00111001000000000000000000000",
		--Instruccion NOPE
		15 => "00111100000000000000000000000",
		--Operations
		16 => "00110011001000000000000000101", -- 5 X
		17 => "00111010001000000000000000010", -- 2 Y
		18 => "00111010001000000000000000001", -- 1 Z
		19 => "00101011001000000000111110100", -- 500 W
		others => "00000000000000000000000000000"
	);
begin
	memoryValue <= TR(conv_integer(direction));
end ArchROM;